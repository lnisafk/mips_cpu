`timescale 1ns / 1ps
module IFU(
    input  clk, rst,
    input  Zero, 
    input  [1:0]  PcSrc,
    input  [31:0] Instr_in,
    input  [31:0] JrAddr,
    output [31:0] JalAddr,
    output [31:0] Instr_out
);
    reg [31:0] ROM[0:31];
    reg [31:0] pc, npc;

    initial pc = 32'h00000000;
    initial $readmemh("code.txt", ROM);
    assign Instr_out = ROM[pc[6:2]];
    assign JalAddr = (PcSrc == 2)?pc+4:0;

    always@(*) begin                        // NPC
        if (PcSrc == 1 && Zero == 1)
            npc <= pc + 4 + (Instr_in[15:0] << 2);
        else if (PcSrc == 2)
            npc <= {pc[31:28], Instr_in[25:0], 2'b00}; 
        else if (PcSrc == 3)
            npc <= JrAddr;
        else
            npc <= pc + 4;
    end

    always@(posedge clk) begin              // PC
        if(rst == 1)
            pc <= 32'h00000000;
        else begin
            pc <= npc;  
            $display("\nPC  -- %h", npc);	
        end
             
    end
	
    /*
    initial begin
        ROM[0] =  32'h3c11cccc;
        ROM[1] =  32'h36723333;
        ROM[2] =  32'h02329821;
        ROM[3] =  32'h0271a023;
        ROM[4] =  32'h12540002;
        ROM[5] =  32'h00000000;
        ROM[6] =  32'hae510004;
        ROM[7] =  32'h8e550004;
        ROM[8] =  32'b000000_00000_00000_00000_00000_000000;
        ROM[9] =  32'b000000_00000_00000_00000_00000_000000;
        ROM[10] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[11] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[12] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[13] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[14] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[15] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[16] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[17] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[18] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[19] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[20] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[21] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[22] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[23] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[24] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[25] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[26] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[27] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[28] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[29] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[30] = 32'b000000_00000_00000_00000_00000_000000;
        ROM[31] = 32'b000000_00000_00000_00000_00000_000000;
    end
    */
endmodule